
module _$_;
    and anon_0 (c_and_d, c, d);
    buf anon_1 (h2, h);
    bufif0 anon_2 (out, in, ctl);
    bufif1 anon_3 (out, in, ctl);
    cmos anon_4 (out, in, nctl, pctl);
    nand anon_5 (d_nand_e, d, e);
    nmos anon_6 (out, in, ctl);
    nor anon_7 (e_nor_f, e, f);
    not anon_8 (a_bar, a);
    notif0 anon_9 (out, in, ctl);
    notif1 anon_10 (out, in, ctl);
    or anon_11 (b_or_c, b, c);
    pmos anon_12 (out, in, ctl);
    pulldown anon_13 (out);
    pullup anon_14 (out);
    rcmos anon_15 (out, in, nctl, pctl);
    rnmos anon_16 (out, in, ctl);
    rpmos anon_17 (out, in, ctl);
    rtran anon_18 (io, io);
    rtranif0 anon_19 (out, in, ctl);
    rtranif1 anon_20 (out, in, ctl);
    tran anon_21 (io, io);
    tranif0 anon_22 (out, in, ctl);
    tranif1 anon_23 (out, in, ctl);
    xnor anon_24 (g_xnor_h, g, h);
    xor anon_25 (f_xor_g, f, g);
endmodule
